`include "base_test.sv"

`include "test_dummy"
//other tests